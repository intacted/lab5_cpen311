module fast_to_slow(
    input clk1,clk2,in,
    output out,
)