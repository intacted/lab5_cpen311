// DE1_SoC_QSYS.v

// Generated using ACDS version 14.1 186 at 2021.04.05.00:40:13

`timescale 1 ps / 1 ps
module DE1_SoC_QSYS (
		output wire [31:0] audio2fifo_0_data_divfrec_export,                  //                  audio2fifo_0_data_divfrec.export
		input  wire        audio2fifo_0_empty_export,                         //                         audio2fifo_0_empty.export
		input  wire        audio2fifo_0_fifo_full_export,                     //                     audio2fifo_0_fifo_full.export
		input  wire [11:0] audio2fifo_0_fifo_used_export,                     //                     audio2fifo_0_fifo_used.export
		output wire [31:0] audio2fifo_0_out_data_audio_export,                //                audio2fifo_0_out_data_audio.export
		output wire        audio2fifo_0_out_pause_export,                     //                     audio2fifo_0_out_pause.export
		output wire        audio2fifo_0_out_stop_export,                      //                      audio2fifo_0_out_stop.export
		output wire        audio2fifo_0_wrclk_export,                         //                         audio2fifo_0_wrclk.export
		output wire        audio2fifo_0_wrreq_export,                         //                         audio2fifo_0_wrreq.export
		output wire        audio_sel_export,                                  //                                  audio_sel.export
		input  wire        clk_clk,                                           //                                        clk.clk
		output wire        clk_25_out_clk,                                    //                                 clk_25_out.clk
		output wire        clk_sdram_clk,                                     //                                  clk_sdram.clk
		output wire [31:0] dds_increment_external_connection_export,          //          dds_increment_external_connection.export
		output wire [31:0] div_freq_export,                                   //                                   div_freq.export
		input  wire [3:0]  key_external_connection_export,                    //                    key_external_connection.export
		input  wire [31:0] keyboard_keys_export,                              //                              keyboard_keys.export
		input  wire        lfsr_clk_interrupt_gen_external_connection_export, // lfsr_clk_interrupt_gen_external_connection.export
		input  wire [31:0] lfsr_val_external_connection_export,               //               lfsr_val_external_connection.export
		output wire [3:0]  modulation_selector_export,                        //                        modulation_selector.export
		input  wire [31:0] mouse_pos_export,                                  //                                  mouse_pos.export
		output wire        pll_locked_export,                                 //                                 pll_locked.export
		input  wire        reset_reset_n,                                     //                                      reset.reset_n
		output wire [12:0] sdram_wire_addr,                                   //                                 sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                     //                                           .ba
		output wire        sdram_wire_cas_n,                                  //                                           .cas_n
		output wire        sdram_wire_cke,                                    //                                           .cke
		output wire        sdram_wire_cs_n,                                   //                                           .cs_n
		inout  wire [15:0] sdram_wire_dq,                                     //                                           .dq
		output wire [1:0]  sdram_wire_dqm,                                    //                                           .dqm
		output wire        sdram_wire_ras_n,                                  //                                           .ras_n
		output wire        sdram_wire_we_n,                                   //                                           .we_n
		output wire [7:0]  signal_selector_export,                            //                            signal_selector.export
		input  wire        vga_alt_vip_itc_0_clocked_video_vid_clk,           //            vga_alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] vga_alt_vip_itc_0_clocked_video_vid_data,          //                                           .vid_data
		output wire        vga_alt_vip_itc_0_clocked_video_underflow,         //                                           .underflow
		output wire        vga_alt_vip_itc_0_clocked_video_vid_datavalid,     //                                           .vid_datavalid
		output wire        vga_alt_vip_itc_0_clocked_video_vid_v_sync,        //                                           .vid_v_sync
		output wire        vga_alt_vip_itc_0_clocked_video_vid_h_sync,        //                                           .vid_h_sync
		output wire        vga_alt_vip_itc_0_clocked_video_vid_f,             //                                           .vid_f
		output wire        vga_alt_vip_itc_0_clocked_video_vid_h,             //                                           .vid_h
		output wire        vga_alt_vip_itc_0_clocked_video_vid_v,             //                                           .vid_v
		output wire        vga_vga_clk_clk                                    //                                vga_vga_clk.clk
	);

	wire         pll_outclk0_clk;                                           // pll:outclk_0 -> [audio:clk_clk, irq_synchronizer:receiver_clk, mm_interconnect_0:pll_outclk0_clk, rst_controller:clk, sdram:clk, vga:nios_clk_clk]
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] vga_to_sdram_readdata;                                     // mm_interconnect_0:vga_to_sdram_readdata -> vga:to_sdram_readdata
	wire         vga_to_sdram_waitrequest;                                  // mm_interconnect_0:vga_to_sdram_waitrequest -> vga:to_sdram_waitrequest
	wire  [31:0] vga_to_sdram_address;                                      // vga:to_sdram_address -> mm_interconnect_0:vga_to_sdram_address
	wire         vga_to_sdram_read;                                         // vga:to_sdram_read -> mm_interconnect_0:vga_to_sdram_read
	wire         vga_to_sdram_readdatavalid;                                // mm_interconnect_0:vga_to_sdram_readdatavalid -> vga:to_sdram_readdatavalid
	wire   [5:0] vga_to_sdram_burstcount;                                   // vga:to_sdram_burstcount -> mm_interconnect_0:vga_to_sdram_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire         mm_interconnect_0_audio_data_fregen_s1_chipselect;         // mm_interconnect_0:audio_data_fregen_s1_chipselect -> audio:data_fregen_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_data_fregen_s1_readdata;           // audio:data_fregen_s1_readdata -> mm_interconnect_0:audio_data_fregen_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_data_fregen_s1_address;            // mm_interconnect_0:audio_data_fregen_s1_address -> audio:data_fregen_s1_address
	wire         mm_interconnect_0_audio_data_fregen_s1_write;              // mm_interconnect_0:audio_data_fregen_s1_write -> audio:data_fregen_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_data_fregen_s1_writedata;          // mm_interconnect_0:audio_data_fregen_s1_writedata -> audio:data_fregen_s1_writedata
	wire  [31:0] mm_interconnect_0_audio_empty_s1_readdata;                 // audio:empty_s1_readdata -> mm_interconnect_0:audio_empty_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_empty_s1_address;                  // mm_interconnect_0:audio_empty_s1_address -> audio:empty_s1_address
	wire  [31:0] mm_interconnect_0_audio_fifo_full_s1_readdata;             // audio:fifo_full_s1_readdata -> mm_interconnect_0:audio_fifo_full_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_fifo_full_s1_address;              // mm_interconnect_0:audio_fifo_full_s1_address -> audio:fifo_full_s1_address
	wire  [31:0] mm_interconnect_0_audio_fifo_used_s1_readdata;             // audio:fifo_used_s1_readdata -> mm_interconnect_0:audio_fifo_used_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_fifo_used_s1_address;              // mm_interconnect_0:audio_fifo_used_s1_address -> audio:fifo_used_s1_address
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire         mm_interconnect_0_audio_out_data_audio_s1_chipselect;      // mm_interconnect_0:audio_out_data_audio_s1_chipselect -> audio:out_data_audio_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_out_data_audio_s1_readdata;        // audio:out_data_audio_s1_readdata -> mm_interconnect_0:audio_out_data_audio_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_out_data_audio_s1_address;         // mm_interconnect_0:audio_out_data_audio_s1_address -> audio:out_data_audio_s1_address
	wire         mm_interconnect_0_audio_out_data_audio_s1_write;           // mm_interconnect_0:audio_out_data_audio_s1_write -> audio:out_data_audio_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_out_data_audio_s1_writedata;       // mm_interconnect_0:audio_out_data_audio_s1_writedata -> audio:out_data_audio_s1_writedata
	wire         mm_interconnect_0_audio_out_pause_s1_chipselect;           // mm_interconnect_0:audio_out_pause_s1_chipselect -> audio:out_pause_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_out_pause_s1_readdata;             // audio:out_pause_s1_readdata -> mm_interconnect_0:audio_out_pause_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_out_pause_s1_address;              // mm_interconnect_0:audio_out_pause_s1_address -> audio:out_pause_s1_address
	wire         mm_interconnect_0_audio_out_pause_s1_write;                // mm_interconnect_0:audio_out_pause_s1_write -> audio:out_pause_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_out_pause_s1_writedata;            // mm_interconnect_0:audio_out_pause_s1_writedata -> audio:out_pause_s1_writedata
	wire         mm_interconnect_0_audio_out_stop_s1_chipselect;            // mm_interconnect_0:audio_out_stop_s1_chipselect -> audio:out_stop_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_out_stop_s1_readdata;              // audio:out_stop_s1_readdata -> mm_interconnect_0:audio_out_stop_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_out_stop_s1_address;               // mm_interconnect_0:audio_out_stop_s1_address -> audio:out_stop_s1_address
	wire         mm_interconnect_0_audio_out_stop_s1_write;                 // mm_interconnect_0:audio_out_stop_s1_write -> audio:out_stop_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_out_stop_s1_writedata;             // mm_interconnect_0:audio_out_stop_s1_writedata -> audio:out_stop_s1_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                       // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                         // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                          // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_write;                            // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                        // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire         mm_interconnect_0_signal_selector_s1_chipselect;           // mm_interconnect_0:signal_selector_s1_chipselect -> signal_selector:chipselect
	wire  [31:0] mm_interconnect_0_signal_selector_s1_readdata;             // signal_selector:readdata -> mm_interconnect_0:signal_selector_s1_readdata
	wire   [1:0] mm_interconnect_0_signal_selector_s1_address;              // mm_interconnect_0:signal_selector_s1_address -> signal_selector:address
	wire         mm_interconnect_0_signal_selector_s1_write;                // mm_interconnect_0:signal_selector_s1_write -> signal_selector:write_n
	wire  [31:0] mm_interconnect_0_signal_selector_s1_writedata;            // mm_interconnect_0:signal_selector_s1_writedata -> signal_selector:writedata
	wire         mm_interconnect_0_modulation_selector_s1_chipselect;       // mm_interconnect_0:modulation_selector_s1_chipselect -> modulation_selector:chipselect
	wire  [31:0] mm_interconnect_0_modulation_selector_s1_readdata;         // modulation_selector:readdata -> mm_interconnect_0:modulation_selector_s1_readdata
	wire   [1:0] mm_interconnect_0_modulation_selector_s1_address;          // mm_interconnect_0:modulation_selector_s1_address -> modulation_selector:address
	wire         mm_interconnect_0_modulation_selector_s1_write;            // mm_interconnect_0:modulation_selector_s1_write -> modulation_selector:write_n
	wire  [31:0] mm_interconnect_0_modulation_selector_s1_writedata;        // mm_interconnect_0:modulation_selector_s1_writedata -> modulation_selector:writedata
	wire  [31:0] mm_interconnect_0_keyboard_keys_s1_readdata;               // keyboard_keys:readdata -> mm_interconnect_0:keyboard_keys_s1_readdata
	wire   [1:0] mm_interconnect_0_keyboard_keys_s1_address;                // mm_interconnect_0:keyboard_keys_s1_address -> keyboard_keys:address
	wire  [31:0] mm_interconnect_0_mouse_pos_s1_readdata;                   // mouse_pos:readdata -> mm_interconnect_0:mouse_pos_s1_readdata
	wire   [1:0] mm_interconnect_0_mouse_pos_s1_address;                    // mm_interconnect_0:mouse_pos_s1_address -> mouse_pos:address
	wire         mm_interconnect_0_div_freq_s1_chipselect;                  // mm_interconnect_0:div_freq_s1_chipselect -> div_freq:chipselect
	wire  [31:0] mm_interconnect_0_div_freq_s1_readdata;                    // div_freq:readdata -> mm_interconnect_0:div_freq_s1_readdata
	wire   [1:0] mm_interconnect_0_div_freq_s1_address;                     // mm_interconnect_0:div_freq_s1_address -> div_freq:address
	wire         mm_interconnect_0_div_freq_s1_write;                       // mm_interconnect_0:div_freq_s1_write -> div_freq:write_n
	wire  [31:0] mm_interconnect_0_div_freq_s1_writedata;                   // mm_interconnect_0:div_freq_s1_writedata -> div_freq:writedata
	wire         mm_interconnect_0_audio_sel_s1_chipselect;                 // mm_interconnect_0:audio_sel_s1_chipselect -> audio_sel:chipselect
	wire  [31:0] mm_interconnect_0_audio_sel_s1_readdata;                   // audio_sel:readdata -> mm_interconnect_0:audio_sel_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_sel_s1_address;                    // mm_interconnect_0:audio_sel_s1_address -> audio_sel:address
	wire         mm_interconnect_0_audio_sel_s1_write;                      // mm_interconnect_0:audio_sel_s1_write -> audio_sel:write_n
	wire  [31:0] mm_interconnect_0_audio_sel_s1_writedata;                  // mm_interconnect_0:audio_sel_s1_writedata -> audio_sel:writedata
	wire         mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect;    // mm_interconnect_0:lfsr_clk_interrupt_gen_s1_chipselect -> lfsr_clk_interrupt_gen:chipselect
	wire  [31:0] mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata;      // lfsr_clk_interrupt_gen:readdata -> mm_interconnect_0:lfsr_clk_interrupt_gen_s1_readdata
	wire   [1:0] mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address;       // mm_interconnect_0:lfsr_clk_interrupt_gen_s1_address -> lfsr_clk_interrupt_gen:address
	wire         mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write;         // mm_interconnect_0:lfsr_clk_interrupt_gen_s1_write -> lfsr_clk_interrupt_gen:write_n
	wire  [31:0] mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata;     // mm_interconnect_0:lfsr_clk_interrupt_gen_s1_writedata -> lfsr_clk_interrupt_gen:writedata
	wire  [31:0] mm_interconnect_0_lfsr_val_s1_readdata;                    // lfsr_val:readdata -> mm_interconnect_0:lfsr_val_s1_readdata
	wire   [1:0] mm_interconnect_0_lfsr_val_s1_address;                     // mm_interconnect_0:lfsr_val_s1_address -> lfsr_val:address
	wire         mm_interconnect_0_dds_increment_s1_chipselect;             // mm_interconnect_0:dds_increment_s1_chipselect -> dds_increment:chipselect
	wire  [31:0] mm_interconnect_0_dds_increment_s1_readdata;               // dds_increment:readdata -> mm_interconnect_0:dds_increment_s1_readdata
	wire   [1:0] mm_interconnect_0_dds_increment_s1_address;                // mm_interconnect_0:dds_increment_s1_address -> dds_increment:address
	wire         mm_interconnect_0_dds_increment_s1_write;                  // mm_interconnect_0:dds_increment_s1_write -> dds_increment:write_n
	wire  [31:0] mm_interconnect_0_dds_increment_s1_writedata;              // mm_interconnect_0:dds_increment_s1_writedata -> dds_increment:writedata
	wire  [31:0] mm_interconnect_0_vga_to_nios_2_datamaster_readdata;       // vga:to_nios_2_datamaster_readdata -> mm_interconnect_0:vga_to_nios_2_datamaster_readdata
	wire   [4:0] mm_interconnect_0_vga_to_nios_2_datamaster_address;        // mm_interconnect_0:vga_to_nios_2_datamaster_address -> vga:to_nios_2_datamaster_address
	wire         mm_interconnect_0_vga_to_nios_2_datamaster_read;           // mm_interconnect_0:vga_to_nios_2_datamaster_read -> vga:to_nios_2_datamaster_read
	wire         mm_interconnect_0_vga_to_nios_2_datamaster_write;          // mm_interconnect_0:vga_to_nios_2_datamaster_write -> vga:to_nios_2_datamaster_write
	wire  [31:0] mm_interconnect_0_vga_to_nios_2_datamaster_writedata;      // mm_interconnect_0:vga_to_nios_2_datamaster_writedata -> vga:to_nios_2_datamaster_writedata
	wire         mm_interconnect_0_audio_wrclk_s1_chipselect;               // mm_interconnect_0:audio_wrclk_s1_chipselect -> audio:wrclk_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_wrclk_s1_readdata;                 // audio:wrclk_s1_readdata -> mm_interconnect_0:audio_wrclk_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_wrclk_s1_address;                  // mm_interconnect_0:audio_wrclk_s1_address -> audio:wrclk_s1_address
	wire         mm_interconnect_0_audio_wrclk_s1_write;                    // mm_interconnect_0:audio_wrclk_s1_write -> audio:wrclk_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_wrclk_s1_writedata;                // mm_interconnect_0:audio_wrclk_s1_writedata -> audio:wrclk_s1_writedata
	wire         mm_interconnect_0_audio_wrreq_s1_chipselect;               // mm_interconnect_0:audio_wrreq_s1_chipselect -> audio:wrreq_s1_chipselect
	wire  [31:0] mm_interconnect_0_audio_wrreq_s1_readdata;                 // audio:wrreq_s1_readdata -> mm_interconnect_0:audio_wrreq_s1_readdata
	wire   [1:0] mm_interconnect_0_audio_wrreq_s1_address;                  // mm_interconnect_0:audio_wrreq_s1_address -> audio:wrreq_s1_address
	wire         mm_interconnect_0_audio_wrreq_s1_write;                    // mm_interconnect_0:audio_wrreq_s1_write -> audio:wrreq_s1_write_n
	wire  [31:0] mm_interconnect_0_audio_wrreq_s1_writedata;                // mm_interconnect_0:audio_wrreq_s1_writedata -> audio:wrreq_s1_writedata
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // key:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // lfsr_clk_interrupt_gen:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // vga:alt_vip_vfr_0_interrupt_sender_irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [audio:reset_reset_n, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset, mm_interconnect_0:vga_nios_clk_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [audio_sel:reset_n, dds_increment:reset_n, div_freq:reset_n, jtag_uart:rst_n, key:reset_n, lfsr_clk_interrupt_gen:reset_n, lfsr_val:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, modulation_selector:reset_n, signal_selector:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                    // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                         // cpu:jtag_debug_module_resetrequest -> rst_controller_002:reset_in1
	wire         rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [keyboard_keys:reset_n, mm_interconnect_0:keyboard_keys_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                        // rst_controller_004:reset_out -> [mm_interconnect_0:mouse_pos_reset_reset_bridge_in_reset_reset, mouse_pos:reset_n]

	DE1_SoC_QSYS_audio audio (
		.clk_clk                      (pll_outclk0_clk),                                      //               clk.clk
		.data_divfrec_export          (audio2fifo_0_data_divfrec_export),                     //      data_divfrec.export
		.data_fregen_s1_address       (mm_interconnect_0_audio_data_fregen_s1_address),       //    data_fregen_s1.address
		.data_fregen_s1_write_n       (~mm_interconnect_0_audio_data_fregen_s1_write),        //                  .write_n
		.data_fregen_s1_writedata     (mm_interconnect_0_audio_data_fregen_s1_writedata),     //                  .writedata
		.data_fregen_s1_chipselect    (mm_interconnect_0_audio_data_fregen_s1_chipselect),    //                  .chipselect
		.data_fregen_s1_readdata      (mm_interconnect_0_audio_data_fregen_s1_readdata),      //                  .readdata
		.empty_export                 (audio2fifo_0_empty_export),                            //             empty.export
		.empty_s1_address             (mm_interconnect_0_audio_empty_s1_address),             //          empty_s1.address
		.empty_s1_readdata            (mm_interconnect_0_audio_empty_s1_readdata),            //                  .readdata
		.fifo_full_export             (audio2fifo_0_fifo_full_export),                        //         fifo_full.export
		.fifo_full_s1_address         (mm_interconnect_0_audio_fifo_full_s1_address),         //      fifo_full_s1.address
		.fifo_full_s1_readdata        (mm_interconnect_0_audio_fifo_full_s1_readdata),        //                  .readdata
		.fifo_used_export             (audio2fifo_0_fifo_used_export),                        //         fifo_used.export
		.fifo_used_s1_address         (mm_interconnect_0_audio_fifo_used_s1_address),         //      fifo_used_s1.address
		.fifo_used_s1_readdata        (mm_interconnect_0_audio_fifo_used_s1_readdata),        //                  .readdata
		.out_data_audio_export        (audio2fifo_0_out_data_audio_export),                   //    out_data_audio.export
		.out_data_audio_s1_address    (mm_interconnect_0_audio_out_data_audio_s1_address),    // out_data_audio_s1.address
		.out_data_audio_s1_write_n    (~mm_interconnect_0_audio_out_data_audio_s1_write),     //                  .write_n
		.out_data_audio_s1_writedata  (mm_interconnect_0_audio_out_data_audio_s1_writedata),  //                  .writedata
		.out_data_audio_s1_chipselect (mm_interconnect_0_audio_out_data_audio_s1_chipselect), //                  .chipselect
		.out_data_audio_s1_readdata   (mm_interconnect_0_audio_out_data_audio_s1_readdata),   //                  .readdata
		.out_pause_export             (audio2fifo_0_out_pause_export),                        //         out_pause.export
		.out_pause_s1_address         (mm_interconnect_0_audio_out_pause_s1_address),         //      out_pause_s1.address
		.out_pause_s1_write_n         (~mm_interconnect_0_audio_out_pause_s1_write),          //                  .write_n
		.out_pause_s1_writedata       (mm_interconnect_0_audio_out_pause_s1_writedata),       //                  .writedata
		.out_pause_s1_chipselect      (mm_interconnect_0_audio_out_pause_s1_chipselect),      //                  .chipselect
		.out_pause_s1_readdata        (mm_interconnect_0_audio_out_pause_s1_readdata),        //                  .readdata
		.out_stop_export              (audio2fifo_0_out_stop_export),                         //          out_stop.export
		.out_stop_s1_address          (mm_interconnect_0_audio_out_stop_s1_address),          //       out_stop_s1.address
		.out_stop_s1_write_n          (~mm_interconnect_0_audio_out_stop_s1_write),           //                  .write_n
		.out_stop_s1_writedata        (mm_interconnect_0_audio_out_stop_s1_writedata),        //                  .writedata
		.out_stop_s1_chipselect       (mm_interconnect_0_audio_out_stop_s1_chipselect),       //                  .chipselect
		.out_stop_s1_readdata         (mm_interconnect_0_audio_out_stop_s1_readdata),         //                  .readdata
		.reset_reset_n                (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.wrclk_export                 (audio2fifo_0_wrclk_export),                            //             wrclk.export
		.wrclk_s1_address             (mm_interconnect_0_audio_wrclk_s1_address),             //          wrclk_s1.address
		.wrclk_s1_write_n             (~mm_interconnect_0_audio_wrclk_s1_write),              //                  .write_n
		.wrclk_s1_writedata           (mm_interconnect_0_audio_wrclk_s1_writedata),           //                  .writedata
		.wrclk_s1_chipselect          (mm_interconnect_0_audio_wrclk_s1_chipselect),          //                  .chipselect
		.wrclk_s1_readdata            (mm_interconnect_0_audio_wrclk_s1_readdata),            //                  .readdata
		.wrreq_export                 (audio2fifo_0_wrreq_export),                            //             wrreq.export
		.wrreq_s1_address             (mm_interconnect_0_audio_wrreq_s1_address),             //          wrreq_s1.address
		.wrreq_s1_write_n             (~mm_interconnect_0_audio_wrreq_s1_write),              //                  .write_n
		.wrreq_s1_writedata           (mm_interconnect_0_audio_wrreq_s1_writedata),           //                  .writedata
		.wrreq_s1_chipselect          (mm_interconnect_0_audio_wrreq_s1_chipselect),          //                  .chipselect
		.wrreq_s1_readdata            (mm_interconnect_0_audio_wrreq_s1_readdata)             //                  .readdata
	);

	DE1_SoC_QSYS_audio_sel audio_sel (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_audio_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_audio_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_audio_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_audio_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_audio_sel_s1_readdata),   //                    .readdata
		.out_port   (audio_sel_export)                           // external_connection.export
	);

	DE1_SoC_QSYS_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE1_SoC_QSYS_dds_increment dds_increment (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_dds_increment_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dds_increment_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dds_increment_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dds_increment_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dds_increment_s1_readdata),   //                    .readdata
		.out_port   (dds_increment_external_connection_export)       // external_connection.export
	);

	DE1_SoC_QSYS_dds_increment div_freq (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_div_freq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_div_freq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_div_freq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_div_freq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_div_freq_s1_readdata),   //                    .readdata
		.out_port   (div_freq_export)                           // external_connection.export
	);

	DE1_SoC_QSYS_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	DE1_SoC_QSYS_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)             //                 irq.irq
	);

	DE1_SoC_QSYS_keyboard_keys keyboard_keys (
		.clk      (clk_25_out_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_keyboard_keys_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keyboard_keys_s1_readdata), //                    .readdata
		.in_port  (keyboard_keys_export)                         // external_connection.export
	);

	DE1_SoC_QSYS_lfsr_clk_interrupt_gen lfsr_clk_interrupt_gen (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata),   //                    .readdata
		.in_port    (lfsr_clk_interrupt_gen_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                                //                 irq.irq
	);

	DE1_SoC_QSYS_lfsr_val lfsr_val (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_lfsr_val_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lfsr_val_s1_readdata), //                    .readdata
		.in_port  (lfsr_val_external_connection_export)     // external_connection.export
	);

	DE1_SoC_QSYS_modulation_selector modulation_selector (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_modulation_selector_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_modulation_selector_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_modulation_selector_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_modulation_selector_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_modulation_selector_s1_readdata),   //                    .readdata
		.out_port   (modulation_selector_export)                           // external_connection.export
	);

	DE1_SoC_QSYS_mouse_pos mouse_pos (
		.clk      (vga_vga_clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_mouse_pos_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_mouse_pos_s1_readdata), //                    .readdata
		.in_port  (mouse_pos_export)                         // external_connection.export
	);

	DE1_SoC_QSYS_pll pll (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_outclk0_clk),   // outclk0.clk
		.outclk_1 (clk_sdram_clk),     // outclk1.clk
		.outclk_2 (clk_25_out_clk),    // outclk2.clk
		.locked   (pll_locked_export)  //  locked.export
	);

	DE1_SoC_QSYS_sdram sdram (
		.clk            (pll_outclk0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	DE1_SoC_QSYS_signal_selector signal_selector (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_signal_selector_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_signal_selector_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_signal_selector_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_signal_selector_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_signal_selector_s1_readdata),   //                    .readdata
		.out_port   (signal_selector_export)                           // external_connection.export
	);

	DE1_SoC_QSYS_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	DE1_SoC_QSYS_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	DE1_SoC_QSYS_vga vga (
		.alt_vip_itc_0_clocked_video_vid_clk       (vga_alt_vip_itc_0_clocked_video_vid_clk),              //    alt_vip_itc_0_clocked_video.vid_clk
		.alt_vip_itc_0_clocked_video_vid_data      (vga_alt_vip_itc_0_clocked_video_vid_data),             //                               .vid_data
		.alt_vip_itc_0_clocked_video_underflow     (vga_alt_vip_itc_0_clocked_video_underflow),            //                               .underflow
		.alt_vip_itc_0_clocked_video_vid_datavalid (vga_alt_vip_itc_0_clocked_video_vid_datavalid),        //                               .vid_datavalid
		.alt_vip_itc_0_clocked_video_vid_v_sync    (vga_alt_vip_itc_0_clocked_video_vid_v_sync),           //                               .vid_v_sync
		.alt_vip_itc_0_clocked_video_vid_h_sync    (vga_alt_vip_itc_0_clocked_video_vid_h_sync),           //                               .vid_h_sync
		.alt_vip_itc_0_clocked_video_vid_f         (vga_alt_vip_itc_0_clocked_video_vid_f),                //                               .vid_f
		.alt_vip_itc_0_clocked_video_vid_h         (vga_alt_vip_itc_0_clocked_video_vid_h),                //                               .vid_h
		.alt_vip_itc_0_clocked_video_vid_v         (vga_alt_vip_itc_0_clocked_video_vid_v),                //                               .vid_v
		.alt_vip_vfr_0_interrupt_sender_irq        (irq_synchronizer_receiver_irq),                        // alt_vip_vfr_0_interrupt_sender.irq
		.clk_50m_clk                               (clk_clk),                                              //                        clk_50m.clk
		.clk_50m_reset_reset_n                     (reset_reset_n),                                        //                  clk_50m_reset.reset_n
		.nios_clk_clk                              (pll_outclk0_clk),                                      //                       nios_clk.clk
		.nios_clk_reset_reset_n                    (reset_reset_n),                                        //                 nios_clk_reset.reset_n
		.to_nios_2_datamaster_address              (mm_interconnect_0_vga_to_nios_2_datamaster_address),   //           to_nios_2_datamaster.address
		.to_nios_2_datamaster_write                (mm_interconnect_0_vga_to_nios_2_datamaster_write),     //                               .write
		.to_nios_2_datamaster_writedata            (mm_interconnect_0_vga_to_nios_2_datamaster_writedata), //                               .writedata
		.to_nios_2_datamaster_read                 (mm_interconnect_0_vga_to_nios_2_datamaster_read),      //                               .read
		.to_nios_2_datamaster_readdata             (mm_interconnect_0_vga_to_nios_2_datamaster_readdata),  //                               .readdata
		.to_sdram_address                          (vga_to_sdram_address),                                 //                       to_sdram.address
		.to_sdram_burstcount                       (vga_to_sdram_burstcount),                              //                               .burstcount
		.to_sdram_readdata                         (vga_to_sdram_readdata),                                //                               .readdata
		.to_sdram_read                             (vga_to_sdram_read),                                    //                               .read
		.to_sdram_readdatavalid                    (vga_to_sdram_readdatavalid),                           //                               .readdatavalid
		.to_sdram_waitrequest                      (vga_to_sdram_waitrequest),                             //                               .waitrequest
		.vga_clk_clk                               (vga_vga_clk_clk)                                       //                        vga_clk.clk
	);

	DE1_SoC_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                  (clk_clk),                                                   //                                clk_50_clk.clk
		.pll_outclk0_clk                                 (pll_outclk0_clk),                                           //                               pll_outclk0.clk
		.pll_outclk2_clk                                 (clk_25_out_clk),                                            //                               pll_outclk2.clk
		.vga_clk_bridge_out_out_clk_1_clk                (vga_vga_clk_clk),                                           //              vga_clk_bridge_out_out_clk_1.clk
		.audio_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                            //         audio_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                        //         cpu_reset_n_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                        //     jtag_uart_reset_reset_bridge_in_reset.reset
		.keyboard_keys_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                        // keyboard_keys_reset_reset_bridge_in_reset.reset
		.mouse_pos_reset_reset_bridge_in_reset_reset     (rst_controller_004_reset_out_reset),                        //     mouse_pos_reset_reset_bridge_in_reset.reset
		.vga_nios_clk_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                            //  vga_nios_clk_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                         (cpu_data_master_address),                                   //                           cpu_data_master.address
		.cpu_data_master_waitrequest                     (cpu_data_master_waitrequest),                               //                                          .waitrequest
		.cpu_data_master_byteenable                      (cpu_data_master_byteenable),                                //                                          .byteenable
		.cpu_data_master_read                            (cpu_data_master_read),                                      //                                          .read
		.cpu_data_master_readdata                        (cpu_data_master_readdata),                                  //                                          .readdata
		.cpu_data_master_readdatavalid                   (cpu_data_master_readdatavalid),                             //                                          .readdatavalid
		.cpu_data_master_write                           (cpu_data_master_write),                                     //                                          .write
		.cpu_data_master_writedata                       (cpu_data_master_writedata),                                 //                                          .writedata
		.cpu_data_master_debugaccess                     (cpu_data_master_debugaccess),                               //                                          .debugaccess
		.cpu_instruction_master_address                  (cpu_instruction_master_address),                            //                    cpu_instruction_master.address
		.cpu_instruction_master_waitrequest              (cpu_instruction_master_waitrequest),                        //                                          .waitrequest
		.cpu_instruction_master_read                     (cpu_instruction_master_read),                               //                                          .read
		.cpu_instruction_master_readdata                 (cpu_instruction_master_readdata),                           //                                          .readdata
		.cpu_instruction_master_readdatavalid            (cpu_instruction_master_readdatavalid),                      //                                          .readdatavalid
		.vga_to_sdram_address                            (vga_to_sdram_address),                                      //                              vga_to_sdram.address
		.vga_to_sdram_waitrequest                        (vga_to_sdram_waitrequest),                                  //                                          .waitrequest
		.vga_to_sdram_burstcount                         (vga_to_sdram_burstcount),                                   //                                          .burstcount
		.vga_to_sdram_read                               (vga_to_sdram_read),                                         //                                          .read
		.vga_to_sdram_readdata                           (vga_to_sdram_readdata),                                     //                                          .readdata
		.vga_to_sdram_readdatavalid                      (vga_to_sdram_readdatavalid),                                //                                          .readdatavalid
		.audio_data_fregen_s1_address                    (mm_interconnect_0_audio_data_fregen_s1_address),            //                      audio_data_fregen_s1.address
		.audio_data_fregen_s1_write                      (mm_interconnect_0_audio_data_fregen_s1_write),              //                                          .write
		.audio_data_fregen_s1_readdata                   (mm_interconnect_0_audio_data_fregen_s1_readdata),           //                                          .readdata
		.audio_data_fregen_s1_writedata                  (mm_interconnect_0_audio_data_fregen_s1_writedata),          //                                          .writedata
		.audio_data_fregen_s1_chipselect                 (mm_interconnect_0_audio_data_fregen_s1_chipselect),         //                                          .chipselect
		.audio_empty_s1_address                          (mm_interconnect_0_audio_empty_s1_address),                  //                            audio_empty_s1.address
		.audio_empty_s1_readdata                         (mm_interconnect_0_audio_empty_s1_readdata),                 //                                          .readdata
		.audio_fifo_full_s1_address                      (mm_interconnect_0_audio_fifo_full_s1_address),              //                        audio_fifo_full_s1.address
		.audio_fifo_full_s1_readdata                     (mm_interconnect_0_audio_fifo_full_s1_readdata),             //                                          .readdata
		.audio_fifo_used_s1_address                      (mm_interconnect_0_audio_fifo_used_s1_address),              //                        audio_fifo_used_s1.address
		.audio_fifo_used_s1_readdata                     (mm_interconnect_0_audio_fifo_used_s1_readdata),             //                                          .readdata
		.audio_out_data_audio_s1_address                 (mm_interconnect_0_audio_out_data_audio_s1_address),         //                   audio_out_data_audio_s1.address
		.audio_out_data_audio_s1_write                   (mm_interconnect_0_audio_out_data_audio_s1_write),           //                                          .write
		.audio_out_data_audio_s1_readdata                (mm_interconnect_0_audio_out_data_audio_s1_readdata),        //                                          .readdata
		.audio_out_data_audio_s1_writedata               (mm_interconnect_0_audio_out_data_audio_s1_writedata),       //                                          .writedata
		.audio_out_data_audio_s1_chipselect              (mm_interconnect_0_audio_out_data_audio_s1_chipselect),      //                                          .chipselect
		.audio_out_pause_s1_address                      (mm_interconnect_0_audio_out_pause_s1_address),              //                        audio_out_pause_s1.address
		.audio_out_pause_s1_write                        (mm_interconnect_0_audio_out_pause_s1_write),                //                                          .write
		.audio_out_pause_s1_readdata                     (mm_interconnect_0_audio_out_pause_s1_readdata),             //                                          .readdata
		.audio_out_pause_s1_writedata                    (mm_interconnect_0_audio_out_pause_s1_writedata),            //                                          .writedata
		.audio_out_pause_s1_chipselect                   (mm_interconnect_0_audio_out_pause_s1_chipselect),           //                                          .chipselect
		.audio_out_stop_s1_address                       (mm_interconnect_0_audio_out_stop_s1_address),               //                         audio_out_stop_s1.address
		.audio_out_stop_s1_write                         (mm_interconnect_0_audio_out_stop_s1_write),                 //                                          .write
		.audio_out_stop_s1_readdata                      (mm_interconnect_0_audio_out_stop_s1_readdata),              //                                          .readdata
		.audio_out_stop_s1_writedata                     (mm_interconnect_0_audio_out_stop_s1_writedata),             //                                          .writedata
		.audio_out_stop_s1_chipselect                    (mm_interconnect_0_audio_out_stop_s1_chipselect),            //                                          .chipselect
		.audio_wrclk_s1_address                          (mm_interconnect_0_audio_wrclk_s1_address),                  //                            audio_wrclk_s1.address
		.audio_wrclk_s1_write                            (mm_interconnect_0_audio_wrclk_s1_write),                    //                                          .write
		.audio_wrclk_s1_readdata                         (mm_interconnect_0_audio_wrclk_s1_readdata),                 //                                          .readdata
		.audio_wrclk_s1_writedata                        (mm_interconnect_0_audio_wrclk_s1_writedata),                //                                          .writedata
		.audio_wrclk_s1_chipselect                       (mm_interconnect_0_audio_wrclk_s1_chipselect),               //                                          .chipselect
		.audio_wrreq_s1_address                          (mm_interconnect_0_audio_wrreq_s1_address),                  //                            audio_wrreq_s1.address
		.audio_wrreq_s1_write                            (mm_interconnect_0_audio_wrreq_s1_write),                    //                                          .write
		.audio_wrreq_s1_readdata                         (mm_interconnect_0_audio_wrreq_s1_readdata),                 //                                          .readdata
		.audio_wrreq_s1_writedata                        (mm_interconnect_0_audio_wrreq_s1_writedata),                //                                          .writedata
		.audio_wrreq_s1_chipselect                       (mm_interconnect_0_audio_wrreq_s1_chipselect),               //                                          .chipselect
		.audio_sel_s1_address                            (mm_interconnect_0_audio_sel_s1_address),                    //                              audio_sel_s1.address
		.audio_sel_s1_write                              (mm_interconnect_0_audio_sel_s1_write),                      //                                          .write
		.audio_sel_s1_readdata                           (mm_interconnect_0_audio_sel_s1_readdata),                   //                                          .readdata
		.audio_sel_s1_writedata                          (mm_interconnect_0_audio_sel_s1_writedata),                  //                                          .writedata
		.audio_sel_s1_chipselect                         (mm_interconnect_0_audio_sel_s1_chipselect),                 //                                          .chipselect
		.cpu_jtag_debug_module_address                   (mm_interconnect_0_cpu_jtag_debug_module_address),           //                     cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                     (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                          .write
		.cpu_jtag_debug_module_read                      (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                          .read
		.cpu_jtag_debug_module_readdata                  (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                          .readdata
		.cpu_jtag_debug_module_writedata                 (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                          .writedata
		.cpu_jtag_debug_module_byteenable                (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                          .byteenable
		.cpu_jtag_debug_module_waitrequest               (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                          .waitrequest
		.cpu_jtag_debug_module_debugaccess               (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                          .debugaccess
		.dds_increment_s1_address                        (mm_interconnect_0_dds_increment_s1_address),                //                          dds_increment_s1.address
		.dds_increment_s1_write                          (mm_interconnect_0_dds_increment_s1_write),                  //                                          .write
		.dds_increment_s1_readdata                       (mm_interconnect_0_dds_increment_s1_readdata),               //                                          .readdata
		.dds_increment_s1_writedata                      (mm_interconnect_0_dds_increment_s1_writedata),              //                                          .writedata
		.dds_increment_s1_chipselect                     (mm_interconnect_0_dds_increment_s1_chipselect),             //                                          .chipselect
		.div_freq_s1_address                             (mm_interconnect_0_div_freq_s1_address),                     //                               div_freq_s1.address
		.div_freq_s1_write                               (mm_interconnect_0_div_freq_s1_write),                       //                                          .write
		.div_freq_s1_readdata                            (mm_interconnect_0_div_freq_s1_readdata),                    //                                          .readdata
		.div_freq_s1_writedata                           (mm_interconnect_0_div_freq_s1_writedata),                   //                                          .writedata
		.div_freq_s1_chipselect                          (mm_interconnect_0_div_freq_s1_chipselect),                  //                                          .chipselect
		.jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //               jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.key_s1_address                                  (mm_interconnect_0_key_s1_address),                          //                                    key_s1.address
		.key_s1_write                                    (mm_interconnect_0_key_s1_write),                            //                                          .write
		.key_s1_readdata                                 (mm_interconnect_0_key_s1_readdata),                         //                                          .readdata
		.key_s1_writedata                                (mm_interconnect_0_key_s1_writedata),                        //                                          .writedata
		.key_s1_chipselect                               (mm_interconnect_0_key_s1_chipselect),                       //                                          .chipselect
		.keyboard_keys_s1_address                        (mm_interconnect_0_keyboard_keys_s1_address),                //                          keyboard_keys_s1.address
		.keyboard_keys_s1_readdata                       (mm_interconnect_0_keyboard_keys_s1_readdata),               //                                          .readdata
		.lfsr_clk_interrupt_gen_s1_address               (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address),       //                 lfsr_clk_interrupt_gen_s1.address
		.lfsr_clk_interrupt_gen_s1_write                 (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write),         //                                          .write
		.lfsr_clk_interrupt_gen_s1_readdata              (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata),      //                                          .readdata
		.lfsr_clk_interrupt_gen_s1_writedata             (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata),     //                                          .writedata
		.lfsr_clk_interrupt_gen_s1_chipselect            (mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect),    //                                          .chipselect
		.lfsr_val_s1_address                             (mm_interconnect_0_lfsr_val_s1_address),                     //                               lfsr_val_s1.address
		.lfsr_val_s1_readdata                            (mm_interconnect_0_lfsr_val_s1_readdata),                    //                                          .readdata
		.modulation_selector_s1_address                  (mm_interconnect_0_modulation_selector_s1_address),          //                    modulation_selector_s1.address
		.modulation_selector_s1_write                    (mm_interconnect_0_modulation_selector_s1_write),            //                                          .write
		.modulation_selector_s1_readdata                 (mm_interconnect_0_modulation_selector_s1_readdata),         //                                          .readdata
		.modulation_selector_s1_writedata                (mm_interconnect_0_modulation_selector_s1_writedata),        //                                          .writedata
		.modulation_selector_s1_chipselect               (mm_interconnect_0_modulation_selector_s1_chipselect),       //                                          .chipselect
		.mouse_pos_s1_address                            (mm_interconnect_0_mouse_pos_s1_address),                    //                              mouse_pos_s1.address
		.mouse_pos_s1_readdata                           (mm_interconnect_0_mouse_pos_s1_readdata),                   //                                          .readdata
		.sdram_s1_address                                (mm_interconnect_0_sdram_s1_address),                        //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_0_sdram_s1_write),                          //                                          .write
		.sdram_s1_read                                   (mm_interconnect_0_sdram_s1_read),                           //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_0_sdram_s1_readdata),                       //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_0_sdram_s1_writedata),                      //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_0_sdram_s1_byteenable),                     //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_0_sdram_s1_waitrequest),                    //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_0_sdram_s1_chipselect),                     //                                          .chipselect
		.signal_selector_s1_address                      (mm_interconnect_0_signal_selector_s1_address),              //                        signal_selector_s1.address
		.signal_selector_s1_write                        (mm_interconnect_0_signal_selector_s1_write),                //                                          .write
		.signal_selector_s1_readdata                     (mm_interconnect_0_signal_selector_s1_readdata),             //                                          .readdata
		.signal_selector_s1_writedata                    (mm_interconnect_0_signal_selector_s1_writedata),            //                                          .writedata
		.signal_selector_s1_chipselect                   (mm_interconnect_0_signal_selector_s1_chipselect),           //                                          .chipselect
		.sysid_qsys_control_slave_address                (mm_interconnect_0_sysid_qsys_control_slave_address),        //                  sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata               (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                          .readdata
		.timer_s1_address                                (mm_interconnect_0_timer_s1_address),                        //                                  timer_s1.address
		.timer_s1_write                                  (mm_interconnect_0_timer_s1_write),                          //                                          .write
		.timer_s1_readdata                               (mm_interconnect_0_timer_s1_readdata),                       //                                          .readdata
		.timer_s1_writedata                              (mm_interconnect_0_timer_s1_writedata),                      //                                          .writedata
		.timer_s1_chipselect                             (mm_interconnect_0_timer_s1_chipselect),                     //                                          .chipselect
		.vga_to_nios_2_datamaster_address                (mm_interconnect_0_vga_to_nios_2_datamaster_address),        //                  vga_to_nios_2_datamaster.address
		.vga_to_nios_2_datamaster_write                  (mm_interconnect_0_vga_to_nios_2_datamaster_write),          //                                          .write
		.vga_to_nios_2_datamaster_read                   (mm_interconnect_0_vga_to_nios_2_datamaster_read),           //                                          .read
		.vga_to_nios_2_datamaster_readdata               (mm_interconnect_0_vga_to_nios_2_datamaster_readdata),       //                                          .readdata
		.vga_to_nios_2_datamaster_writedata              (mm_interconnect_0_vga_to_nios_2_datamaster_writedata)       //                                          .writedata
	);

	DE1_SoC_QSYS_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_outclk0_clk),                    //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_25_out_clk),                     //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (vga_vga_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
