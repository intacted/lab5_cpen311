// DE1_SoC_QSYS_tb.v

// Generated using ACDS version 14.1 186 at 2021.04.04.17:55:37

`timescale 1 ps / 1 ps
module DE1_SoC_QSYS_tb (
	);

	wire         de1_soc_qsys_inst_clk_bfm_clk_clk;                                               // DE1_SoC_QSYS_inst_clk_bfm:clk -> [DE1_SoC_QSYS_inst:clk_clk, DE1_SoC_QSYS_inst_reset_bfm:clk]
	wire         sdram_my_partner_clk_bfm_clk_clk;                                                // sdram_my_partner_clk_bfm:clk -> sdram_my_partner:clk
	wire  [31:0] de1_soc_qsys_inst_audio2fifo_0_data_divfrec_export;                              // DE1_SoC_QSYS_inst:audio2fifo_0_data_divfrec_export -> DE1_SoC_QSYS_inst_audio2fifo_0_data_divfrec_bfm:sig_export
	wire   [0:0] de1_soc_qsys_inst_audio2fifo_0_empty_bfm_conduit_export;                         // DE1_SoC_QSYS_inst_audio2fifo_0_empty_bfm:sig_export -> DE1_SoC_QSYS_inst:audio2fifo_0_empty_export
	wire   [0:0] de1_soc_qsys_inst_audio2fifo_0_fifo_full_bfm_conduit_export;                     // DE1_SoC_QSYS_inst_audio2fifo_0_fifo_full_bfm:sig_export -> DE1_SoC_QSYS_inst:audio2fifo_0_fifo_full_export
	wire  [11:0] de1_soc_qsys_inst_audio2fifo_0_fifo_used_bfm_conduit_export;                     // DE1_SoC_QSYS_inst_audio2fifo_0_fifo_used_bfm:sig_export -> DE1_SoC_QSYS_inst:audio2fifo_0_fifo_used_export
	wire  [31:0] de1_soc_qsys_inst_audio2fifo_0_out_data_audio_export;                            // DE1_SoC_QSYS_inst:audio2fifo_0_out_data_audio_export -> DE1_SoC_QSYS_inst_audio2fifo_0_out_data_audio_bfm:sig_export
	wire         de1_soc_qsys_inst_audio2fifo_0_out_pause_export;                                 // DE1_SoC_QSYS_inst:audio2fifo_0_out_pause_export -> DE1_SoC_QSYS_inst_audio2fifo_0_out_pause_bfm:sig_export
	wire         de1_soc_qsys_inst_audio2fifo_0_out_stop_export;                                  // DE1_SoC_QSYS_inst:audio2fifo_0_out_stop_export -> DE1_SoC_QSYS_inst_audio2fifo_0_out_stop_bfm:sig_export
	wire         de1_soc_qsys_inst_audio2fifo_0_wrclk_export;                                     // DE1_SoC_QSYS_inst:audio2fifo_0_wrclk_export -> DE1_SoC_QSYS_inst_audio2fifo_0_wrclk_bfm:sig_export
	wire         de1_soc_qsys_inst_audio2fifo_0_wrreq_export;                                     // DE1_SoC_QSYS_inst:audio2fifo_0_wrreq_export -> DE1_SoC_QSYS_inst_audio2fifo_0_wrreq_bfm:sig_export
	wire         de1_soc_qsys_inst_audio_sel_export;                                              // DE1_SoC_QSYS_inst:audio_sel_export -> DE1_SoC_QSYS_inst_audio_sel_bfm:sig_export
	wire  [31:0] de1_soc_qsys_inst_dds_increment_external_connection_export;                      // DE1_SoC_QSYS_inst:dds_increment_external_connection_export -> DE1_SoC_QSYS_inst_dds_increment_external_connection_bfm:sig_export
	wire  [31:0] de1_soc_qsys_inst_div_freq_export;                                               // DE1_SoC_QSYS_inst:div_freq_export -> DE1_SoC_QSYS_inst_div_freq_bfm:sig_export
	wire   [3:0] de1_soc_qsys_inst_key_external_connection_bfm_conduit_export;                    // DE1_SoC_QSYS_inst_key_external_connection_bfm:sig_export -> DE1_SoC_QSYS_inst:key_external_connection_export
	wire  [31:0] de1_soc_qsys_inst_keyboard_keys_bfm_conduit_export;                              // DE1_SoC_QSYS_inst_keyboard_keys_bfm:sig_export -> DE1_SoC_QSYS_inst:keyboard_keys_export
	wire   [0:0] de1_soc_qsys_inst_lfsr_clk_interrupt_gen_external_connection_bfm_conduit_export; // DE1_SoC_QSYS_inst_lfsr_clk_interrupt_gen_external_connection_bfm:sig_export -> DE1_SoC_QSYS_inst:lfsr_clk_interrupt_gen_external_connection_export
	wire  [31:0] de1_soc_qsys_inst_lfsr_val_external_connection_bfm_conduit_export;               // DE1_SoC_QSYS_inst_lfsr_val_external_connection_bfm:sig_export -> DE1_SoC_QSYS_inst:lfsr_val_external_connection_export
	wire   [3:0] de1_soc_qsys_inst_modulation_selector_export;                                    // DE1_SoC_QSYS_inst:modulation_selector_export -> DE1_SoC_QSYS_inst_modulation_selector_bfm:sig_export
	wire  [31:0] de1_soc_qsys_inst_mouse_pos_bfm_conduit_export;                                  // DE1_SoC_QSYS_inst_mouse_pos_bfm:sig_export -> DE1_SoC_QSYS_inst:mouse_pos_export
	wire         de1_soc_qsys_inst_pll_locked_export;                                             // DE1_SoC_QSYS_inst:pll_locked_export -> DE1_SoC_QSYS_inst_pll_locked_bfm:sig_export
	wire         de1_soc_qsys_inst_sdram_wire_cs_n;                                               // DE1_SoC_QSYS_inst:sdram_wire_cs_n -> sdram_my_partner:zs_cs_n
	wire   [1:0] de1_soc_qsys_inst_sdram_wire_dqm;                                                // DE1_SoC_QSYS_inst:sdram_wire_dqm -> sdram_my_partner:zs_dqm
	wire         de1_soc_qsys_inst_sdram_wire_cas_n;                                              // DE1_SoC_QSYS_inst:sdram_wire_cas_n -> sdram_my_partner:zs_cas_n
	wire         de1_soc_qsys_inst_sdram_wire_ras_n;                                              // DE1_SoC_QSYS_inst:sdram_wire_ras_n -> sdram_my_partner:zs_ras_n
	wire         de1_soc_qsys_inst_sdram_wire_we_n;                                               // DE1_SoC_QSYS_inst:sdram_wire_we_n -> sdram_my_partner:zs_we_n
	wire  [12:0] de1_soc_qsys_inst_sdram_wire_addr;                                               // DE1_SoC_QSYS_inst:sdram_wire_addr -> sdram_my_partner:zs_addr
	wire         de1_soc_qsys_inst_sdram_wire_cke;                                                // DE1_SoC_QSYS_inst:sdram_wire_cke -> sdram_my_partner:zs_cke
	wire  [15:0] de1_soc_qsys_inst_sdram_wire_dq;                                                 // [] -> [DE1_SoC_QSYS_inst:sdram_wire_dq, sdram_my_partner:zs_dq]
	wire   [1:0] de1_soc_qsys_inst_sdram_wire_ba;                                                 // DE1_SoC_QSYS_inst:sdram_wire_ba -> sdram_my_partner:zs_ba
	wire   [7:0] de1_soc_qsys_inst_signal_selector_export;                                        // DE1_SoC_QSYS_inst:signal_selector_export -> DE1_SoC_QSYS_inst_signal_selector_bfm:sig_export
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_underflow;                     // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_underflow -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_underflow
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_f;                         // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_f -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_f
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v;                         // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_v -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_v
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h_sync;                    // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_h_sync -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_h_sync
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h;                         // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_h -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_h
	wire   [0:0] de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk;           // DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_clk -> DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_clk
	wire  [23:0] de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_data;                      // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_data -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_data
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_datavalid;                 // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_datavalid -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_datavalid
	wire         de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v_sync;                    // DE1_SoC_QSYS_inst:vga_alt_vip_itc_0_clocked_video_vid_v_sync -> DE1_SoC_QSYS_inst_vga_alt_vip_itc_0_clocked_video_bfm:sig_vid_v_sync
	wire         de1_soc_qsys_inst_reset_bfm_reset_reset;                                         // DE1_SoC_QSYS_inst_reset_bfm:reset -> DE1_SoC_QSYS_inst:reset_reset_n

	DE1_SoC_QSYS de1_soc_qsys_inst (
		.audio2fifo_0_data_divfrec_export                  (de1_soc_qsys_inst_audio2fifo_0_data_divfrec_export),                              //                  audio2fifo_0_data_divfrec.export
		.audio2fifo_0_empty_export                         (de1_soc_qsys_inst_audio2fifo_0_empty_bfm_conduit_export),                         //                         audio2fifo_0_empty.export
		.audio2fifo_0_fifo_full_export                     (de1_soc_qsys_inst_audio2fifo_0_fifo_full_bfm_conduit_export),                     //                     audio2fifo_0_fifo_full.export
		.audio2fifo_0_fifo_used_export                     (de1_soc_qsys_inst_audio2fifo_0_fifo_used_bfm_conduit_export),                     //                     audio2fifo_0_fifo_used.export
		.audio2fifo_0_out_data_audio_export                (de1_soc_qsys_inst_audio2fifo_0_out_data_audio_export),                            //                audio2fifo_0_out_data_audio.export
		.audio2fifo_0_out_pause_export                     (de1_soc_qsys_inst_audio2fifo_0_out_pause_export),                                 //                     audio2fifo_0_out_pause.export
		.audio2fifo_0_out_stop_export                      (de1_soc_qsys_inst_audio2fifo_0_out_stop_export),                                  //                      audio2fifo_0_out_stop.export
		.audio2fifo_0_wrclk_export                         (de1_soc_qsys_inst_audio2fifo_0_wrclk_export),                                     //                         audio2fifo_0_wrclk.export
		.audio2fifo_0_wrreq_export                         (de1_soc_qsys_inst_audio2fifo_0_wrreq_export),                                     //                         audio2fifo_0_wrreq.export
		.audio_sel_export                                  (de1_soc_qsys_inst_audio_sel_export),                                              //                                  audio_sel.export
		.clk_clk                                           (de1_soc_qsys_inst_clk_bfm_clk_clk),                                               //                                        clk.clk
		.clk_25_out_clk                                    (),                                                                                //                                 clk_25_out.clk
		.clk_sdram_clk                                     (),                                                                                //                                  clk_sdram.clk
		.dds_increment_external_connection_export          (de1_soc_qsys_inst_dds_increment_external_connection_export),                      //          dds_increment_external_connection.export
		.div_freq_export                                   (de1_soc_qsys_inst_div_freq_export),                                               //                                   div_freq.export
		.key_external_connection_export                    (de1_soc_qsys_inst_key_external_connection_bfm_conduit_export),                    //                    key_external_connection.export
		.keyboard_keys_export                              (de1_soc_qsys_inst_keyboard_keys_bfm_conduit_export),                              //                              keyboard_keys.export
		.lfsr_clk_interrupt_gen_external_connection_export (de1_soc_qsys_inst_lfsr_clk_interrupt_gen_external_connection_bfm_conduit_export), // lfsr_clk_interrupt_gen_external_connection.export
		.lfsr_val_external_connection_export               (de1_soc_qsys_inst_lfsr_val_external_connection_bfm_conduit_export),               //               lfsr_val_external_connection.export
		.modulation_selector_export                        (de1_soc_qsys_inst_modulation_selector_export),                                    //                        modulation_selector.export
		.mouse_pos_export                                  (de1_soc_qsys_inst_mouse_pos_bfm_conduit_export),                                  //                                  mouse_pos.export
		.pll_locked_export                                 (de1_soc_qsys_inst_pll_locked_export),                                             //                                 pll_locked.export
		.reset_reset_n                                     (de1_soc_qsys_inst_reset_bfm_reset_reset),                                         //                                      reset.reset_n
		.sdram_wire_addr                                   (de1_soc_qsys_inst_sdram_wire_addr),                                               //                                 sdram_wire.addr
		.sdram_wire_ba                                     (de1_soc_qsys_inst_sdram_wire_ba),                                                 //                                           .ba
		.sdram_wire_cas_n                                  (de1_soc_qsys_inst_sdram_wire_cas_n),                                              //                                           .cas_n
		.sdram_wire_cke                                    (de1_soc_qsys_inst_sdram_wire_cke),                                                //                                           .cke
		.sdram_wire_cs_n                                   (de1_soc_qsys_inst_sdram_wire_cs_n),                                               //                                           .cs_n
		.sdram_wire_dq                                     (de1_soc_qsys_inst_sdram_wire_dq),                                                 //                                           .dq
		.sdram_wire_dqm                                    (de1_soc_qsys_inst_sdram_wire_dqm),                                                //                                           .dqm
		.sdram_wire_ras_n                                  (de1_soc_qsys_inst_sdram_wire_ras_n),                                              //                                           .ras_n
		.sdram_wire_we_n                                   (de1_soc_qsys_inst_sdram_wire_we_n),                                               //                                           .we_n
		.signal_selector_export                            (de1_soc_qsys_inst_signal_selector_export),                                        //                            signal_selector.export
		.vga_alt_vip_itc_0_clocked_video_vid_clk           (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk),           //            vga_alt_vip_itc_0_clocked_video.vid_clk
		.vga_alt_vip_itc_0_clocked_video_vid_data          (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_data),                      //                                           .vid_data
		.vga_alt_vip_itc_0_clocked_video_underflow         (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_underflow),                     //                                           .underflow
		.vga_alt_vip_itc_0_clocked_video_vid_datavalid     (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_datavalid),                 //                                           .vid_datavalid
		.vga_alt_vip_itc_0_clocked_video_vid_v_sync        (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v_sync),                    //                                           .vid_v_sync
		.vga_alt_vip_itc_0_clocked_video_vid_h_sync        (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h_sync),                    //                                           .vid_h_sync
		.vga_alt_vip_itc_0_clocked_video_vid_f             (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_f),                         //                                           .vid_f
		.vga_alt_vip_itc_0_clocked_video_vid_h             (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h),                         //                                           .vid_h
		.vga_alt_vip_itc_0_clocked_video_vid_v             (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v),                         //                                           .vid_v
		.vga_vga_clk_clk                                   ()                                                                                 //                                vga_vga_clk.clk
	);

	altera_conduit_bfm de1_soc_qsys_inst_audio2fifo_0_data_divfrec_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_data_divfrec_export)  // conduit.export
	);

	altera_conduit_bfm_0002 de1_soc_qsys_inst_audio2fifo_0_empty_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_empty_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 de1_soc_qsys_inst_audio2fifo_0_fifo_full_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_fifo_full_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 de1_soc_qsys_inst_audio2fifo_0_fifo_used_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_fifo_used_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm de1_soc_qsys_inst_audio2fifo_0_out_data_audio_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_out_data_audio_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_audio2fifo_0_out_pause_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_out_pause_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_audio2fifo_0_out_stop_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_out_stop_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_audio2fifo_0_wrclk_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_wrclk_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_audio2fifo_0_wrreq_bfm (
		.sig_export (de1_soc_qsys_inst_audio2fifo_0_wrreq_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_audio_sel_bfm (
		.sig_export (de1_soc_qsys_inst_audio_sel_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) de1_soc_qsys_inst_clk_bfm (
		.clk (de1_soc_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm de1_soc_qsys_inst_dds_increment_external_connection_bfm (
		.sig_export (de1_soc_qsys_inst_dds_increment_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm de1_soc_qsys_inst_div_freq_bfm (
		.sig_export (de1_soc_qsys_inst_div_freq_export)  // conduit.export
	);

	altera_conduit_bfm_0005 de1_soc_qsys_inst_key_external_connection_bfm (
		.sig_export (de1_soc_qsys_inst_key_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0006 de1_soc_qsys_inst_keyboard_keys_bfm (
		.sig_export (de1_soc_qsys_inst_keyboard_keys_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 de1_soc_qsys_inst_lfsr_clk_interrupt_gen_external_connection_bfm (
		.sig_export (de1_soc_qsys_inst_lfsr_clk_interrupt_gen_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0006 de1_soc_qsys_inst_lfsr_val_external_connection_bfm (
		.sig_export (de1_soc_qsys_inst_lfsr_val_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0007 de1_soc_qsys_inst_modulation_selector_bfm (
		.sig_export (de1_soc_qsys_inst_modulation_selector_export)  // conduit.export
	);

	altera_conduit_bfm_0006 de1_soc_qsys_inst_mouse_pos_bfm (
		.sig_export (de1_soc_qsys_inst_mouse_pos_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de1_soc_qsys_inst_pll_locked_bfm (
		.sig_export (de1_soc_qsys_inst_pll_locked_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) de1_soc_qsys_inst_reset_bfm (
		.reset (de1_soc_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (de1_soc_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0008 de1_soc_qsys_inst_signal_selector_bfm (
		.sig_export (de1_soc_qsys_inst_signal_selector_export)  // conduit.export
	);

	altera_conduit_bfm_0009 de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_bfm (
		.sig_vid_clk       (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk), // conduit.vid_clk
		.sig_vid_data      (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_data),            //        .vid_data
		.sig_underflow     (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_underflow),           //        .underflow
		.sig_vid_datavalid (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_datavalid),       //        .vid_datavalid
		.sig_vid_v_sync    (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v_sync),          //        .vid_v_sync
		.sig_vid_h_sync    (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h_sync),          //        .vid_h_sync
		.sig_vid_f         (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_f),               //        .vid_f
		.sig_vid_h         (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_h),               //        .vid_h
		.sig_vid_v         (de1_soc_qsys_inst_vga_alt_vip_itc_0_clocked_video_vid_v)                //        .vid_v
	);

	altera_sdram_partner_module sdram_my_partner (
		.clk      (sdram_my_partner_clk_bfm_clk_clk),   //     clk.clk
		.zs_dq    (de1_soc_qsys_inst_sdram_wire_dq),    // conduit.dq
		.zs_addr  (de1_soc_qsys_inst_sdram_wire_addr),  //        .addr
		.zs_ba    (de1_soc_qsys_inst_sdram_wire_ba),    //        .ba
		.zs_cas_n (de1_soc_qsys_inst_sdram_wire_cas_n), //        .cas_n
		.zs_cke   (de1_soc_qsys_inst_sdram_wire_cke),   //        .cke
		.zs_cs_n  (de1_soc_qsys_inst_sdram_wire_cs_n),  //        .cs_n
		.zs_dqm   (de1_soc_qsys_inst_sdram_wire_dqm),   //        .dqm
		.zs_ras_n (de1_soc_qsys_inst_sdram_wire_ras_n), //        .ras_n
		.zs_we_n  (de1_soc_qsys_inst_sdram_wire_we_n)   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (142857142),
		.CLOCK_UNIT (1)
	) sdram_my_partner_clk_bfm (
		.clk (sdram_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
